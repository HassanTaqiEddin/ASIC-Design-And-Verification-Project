`ifndef TB_PKG
`define TB_PKG
`include "uvm_macros.svh"
package tb_pkg;
  import uvm_pkg::*;
  
  `include "uvm_macros.svh"
  
  `include "sequence_item.svh"
  `include "sequence.svh"
  `include "sequencer.svh"
  `include "driver.svh"
  `include "monitor.svh"
  `include "scoreboard.svh"
  `include "subscriber.svh"

  `include "agent.svh"
  `include "env.svh"
  `include "test.svh"

endpackage
`endif 
